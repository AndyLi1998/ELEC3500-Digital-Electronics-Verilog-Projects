`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/19/2021 06:25:11 PM
// Design Name: 
// Module Name: lab121
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module lab121(
    input  in0,
    input  in1,
    input  in2,
    input  in3,
    input  in4,
    input  in5,
    input  in6,
    input  in7,
    output out0,
    output out1,
    output out2,
    output out3,
    output out4,
    output out5,
    output out6,
    output out7
    );
    assign out0 = in0;
    assign out1 = in1;
    assign out2 = in2;
    assign out3 = in3;
    assign out4 = in4;
    assign out5 = in5;
    assign out6 = in6;
    assign out7 = in7;
    
endmodule
